// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : Demo01_gen_verilog
// Git hash  : cda2b4527b541defe03b38e53cc3a5260a403089

`timescale 1ns/1ps

module Demo01_gen_verilog (
);



endmodule
