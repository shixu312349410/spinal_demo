// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : Demo04_USint
// Git hash  : 0d5be50c9a8de7ab624975a7e716d258d0b3947c

`timescale 1ns/1ps

module Demo04_USint (
);

  wire       [2:0]    e;
  wire       [3:0]    f;

  assign e = 3'b111;
  assign f = 4'b0111;

endmodule
